-- ============================================================================
-- Grupo de Investigacion en Robotica y Automatizacion Industrial GIRA
-- DescripciÃ³n: 	Memoria con valores constantes de inicializaciÃ³n
-- Autor: 			Wilson Javier PÃ©rez HolguÃ­n
--						Luis Ariel Mesa
--	Fecha:			02-04-2024
-- Estado:			Funcionamiento OK
-- ============================================================================


library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 

entity Memoria_Imagen is

	generic (
		data_width  : natural := 8; 
	   addr_length : natural := 10	-- 1024 pos mem
		); 
	
	port ( 
		clk      :  in std_logic;
--		rst : in std_logic;
		address  :  in std_logic_vector(addr_length-1 downto 0); 
		data_out :  out std_logic_vector(data_width-1  downto 0) 
		);
		
end Memoria_Imagen;


architecture synth of Memoria_Imagen is

	constant mem_size : natural := 2**addr_length; 	
	type mem_type is array (0 to mem_size-1) of std_logic_vector (data_width-1 downto 0); 

constant mem : mem_type := (
		x"02", x"02", x"03", x"03", x"02", x"02", x"01", x"01", x"00", x"06", x"01", x"00", x"02", x"01", x"00", x"02", x"07", x"01", x"00", x"00", x"09", x"02", x"00", x"07", x"04", x"03", x"02", x"01", x"00", x"00", x"00", x"00",
		x"03", x"02", x"01", x"00", x"00", x"02", x"04", x"05", x"07", x"00", x"00", x"07", x"06", x"00", x"00", x"06", x"00", x"08", x"0D", x"08", x"04", x"04", x"03", x"01", x"04", x"03", x"02", x"01", x"00", x"00", x"00", x"00",
		x"04", x"02", x"00", x"00", x"00", x"02", x"05", x"08", x"0A", x"01", x"04", x"0A", x"04", x"03", x"07", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"03", x"04", x"03", x"02", x"01", x"00", x"00", x"00", x"00",
		x"04", x"03", x"02", x"01", x"01", x"02", x"04", x"05", x"03", x"00", x"01", x"00", x"00", x"03", x"0A", x"00", x"13", x"00", x"00", x"07", x"04", x"02", x"03", x"00", x"04", x"03", x"02", x"01", x"00", x"00", x"00", x"00",
		x"03", x"04", x"05", x"05", x"05", x"03", x"01", x"00", x"07", x"04", x"03", x"02", x"01", x"05", x"09", x"05", x"00", x"00", x"02", x"02", x"01", x"06", x"07", x"00", x"04", x"03", x"02", x"01", x"00", x"00", x"00", x"00",
		x"01", x"03", x"06", x"07", x"07", x"04", x"01", x"00", x"02", x"0B", x"16", x"25", x"2B", x"18", x"14", x"2B", x"32", x"50", x"43", x"16", x"04", x"09", x"09", x"07", x"04", x"03", x"02", x"01", x"00", x"00", x"00", x"00",
		x"00", x"01", x"03", x"05", x"06", x"06", x"05", x"05", x"05", x"46", x"6A", x"75", x"83", x"74", x"69", x"83", x"C6", x"DE", x"BF", x"88", x"65", x"30", x"01", x"00", x"04", x"03", x"02", x"01", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"02", x"05", x"07", x"09", x"0A", x"37", x"B7", x"F0", x"E7", x"FB", x"FF", x"F8", x"FF", x"F5", x"FF", x"F3", x"F2", x"E0", x"70", x"05", x"00", x"04", x"03", x"02", x"01", x"00", x"00", x"00", x"00",
		x"06", x"03", x"03", x"05", x"04", x"04", x"09", x"10", x"9C", x"E2", x"FF", x"FF", x"F0", x"FF", x"F9", x"F8", x"FE", x"FC", x"F6", x"FF", x"F8", x"9A", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03",
		x"06", x"03", x"02", x"04", x"04", x"03", x"07", x"0E", x"A3", x"F4", x"F9", x"FF", x"F5", x"F8", x"FB", x"F6", x"FF", x"FF", x"F4", x"F0", x"EF", x"A4", x"08", x"00", x"03", x"04", x"04", x"02", x"00", x"00", x"00", x"02",
		x"05", x"02", x"02", x"03", x"02", x"01", x"04", x"0A", x"74", x"EB", x"F1", x"FE", x"FF", x"FD", x"FF", x"FF", x"F2", x"FF", x"FF", x"F2", x"F4", x"AF", x"04", x"00", x"08", x"08", x"08", x"05", x"01", x"00", x"00", x"01",
		x"04", x"01", x"01", x"03", x"01", x"00", x"02", x"07", x"34", x"C8", x"F7", x"FC", x"E6", x"C8", x"AD", x"B1", x"E8", x"FB", x"FF", x"F8", x"F5", x"AA", x"00", x"0B", x"08", x"09", x"08", x"05", x"01", x"00", x"00", x"01",
		x"03", x"00", x"01", x"02", x"01", x"00", x"01", x"06", x"0B", x"7E", x"D2", x"D7", x"A8", x"6F", x"41", x"86", x"F6", x"F8", x"FB", x"F6", x"EF", x"9D", x"01", x"13", x"05", x"05", x"05", x"03", x"00", x"00", x"00", x"02",
		x"01", x"00", x"00", x"03", x"02", x"00", x"01", x"06", x"00", x"23", x"5F", x"69", x"3F", x"1F", x"27", x"BC", x"FF", x"FA", x"F4", x"FF", x"ED", x"90", x"06", x"05", x"01", x"02", x"03", x"01", x"00", x"00", x"01", x"03",
		x"00", x"00", x"00", x"03", x"03", x"00", x"02", x"07", x"02", x"00", x"08", x"0A", x"00", x"0C", x"4E", x"DF", x"F7", x"FF", x"F6", x"F7", x"C1", x"61", x"04", x"00", x"02", x"03", x"03", x"01", x"00", x"00", x"00", x"02",
		x"00", x"00", x"00", x"04", x"03", x"01", x"03", x"08", x"00", x"0D", x"06", x"0E", x"17", x"56", x"A8", x"F9", x"F2", x"FF", x"F0", x"D2", x"74", x"1F", x"00", x"0C", x"04", x"04", x"04", x"02", x"00", x"00", x"00", x"02",
		x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"05", x"08", x"01", x"00", x"5C", x"D9", x"F6", x"FE", x"F9", x"F9", x"F4", x"6A", x"0E", x"01", x"01", x"07", x"0F", x"03", x"00", x"02", x"03", x"00", x"00", x"03",
		x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"00", x"0E", x"07", x"08", x"67", x"DE", x"FF", x"F5", x"FF", x"DE", x"BE", x"49", x"09", x"08", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"03",
		x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"00", x"07", x"02", x"30", x"95", x"EA", x"FF", x"F3", x"EF", x"72", x"3C", x"08", x"00", x"05", x"09", x"00", x"07", x"0A", x"08", x"01", x"00", x"02", x"02", x"00",
		x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"04", x"01", x"0D", x"74", x"D6", x"F7", x"FF", x"F5", x"EF", x"41", x"02", x"03", x"08", x"00", x"0B", x"0D", x"01", x"00", x"00", x"00", x"00", x"02", x"03", x"03",
		x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"03", x"1B", x"4E", x"BB", x"FA", x"F8", x"FD", x"EE", x"B8", x"27", x"00", x"07", x"08", x"00", x"05", x"00", x"0A", x"00", x"00", x"07", x"0A", x"02", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"48", x"A8", x"EB", x"F8", x"F5", x"F6", x"E1", x"55", x"10", x"04", x"02", x"05", x"09", x"1D", x"06", x"0F", x"0C", x"0B", x"0C", x"07", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5A", x"D3", x"FB", x"F3", x"FC", x"F4", x"DF", x"45", x"25", x"1E", x"15", x"20", x"2E", x"51", x"45", x"4D", x"53", x"41", x"18", x"00", x"00", x"05", x"08",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"4F", x"CE", x"FB", x"FA", x"FF", x"F6", x"E7", x"B3", x"8F", x"83", x"8A", x"A6", x"B6", x"EE", x"FF", x"F9", x"FB", x"C2", x"56", x"09", x"00", x"04", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"37", x"BA", x"FF", x"F7", x"ED", x"F4", x"F8", x"F9", x"F0", x"EE", x"EB", x"E5", x"EE", x"FC", x"FE", x"F9", x"FF", x"C9", x"54", x"00", x"00", x"05", x"04",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"1F", x"86", x"DD", x"FB", x"FF", x"FE", x"F5", x"FD", x"FC", x"FE", x"FE", x"FD", x"FF", x"F3", x"D3", x"90", x"7A", x"48", x"13", x"00", x"09", x"07", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"05", x"42", x"8E", x"D2", x"F9", x"F6", x"F9", x"FB", x"FB", x"FC", x"F5", x"EF", x"E2", x"AF", x"6F", x"2B", x"17", x"02", x"00", x"00", x"05", x"02", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"14", x"36", x"70", x"9A", x"AB", x"CF", x"AD", x"A9", x"A8", x"A4", x"97", x"7F", x"4B", x"0F", x"06", x"05", x"06", x"07", x"01", x"00", x"00", x"06",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"04", x"04", x"01", x"19", x"2D", x"39", x"66", x"33", x"2A", x"30", x"38", x"30", x"21", x"0D", x"00", x"01", x"02", x"00", x"00", x"00", x"04", x"02", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"03", x"00", x"05", x"05", x"00", x"13", x"04", x"00", x"00", x"09", x"02", x"00", x"00", x"06", x"00", x"04", x"02", x"00", x"00", x"05", x"06", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"02", x"09", x"08", x"00", x"02", x"0C", x"05", x"07", x"08", x"00", x"00", x"04", x"04", x"00", x"08", x"0B", x"05", x"00", x"00", x"03", x"06",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"05", x"00", x"06", x"00", x"00", x"03", x"00", x"09", x"00", x"00", x"04", x"02", x"00", x"06", x"07", x"00", x"03", x"00", x"00", x"03", x"04", x"00", x"00", x"00"
	);

	
begin 

	rom : process (clk) 
	begin
	   
----	   if (rising_edge(Clk)) then
--		  if rst = '1' then
--				-- Reset the counter to 0
--				data_out <= ((others=> '0'));
--		  end if;
	   
		if rising_edge(clk) then 
			data_out <= mem(to_integer(unsigned(address))); 
		end if; 
	end process rom; 

end architecture synth;